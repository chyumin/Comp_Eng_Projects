library verilog;
use verilog.vl_types.all;
entity multiplier_seq_vlg_vec_tst is
end multiplier_seq_vlg_vec_tst;
