LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY reg_pp_4bits IS
	PORT (d    :  IN std_logic_vector(3 DOWNTO 0);
			clk  :  IN std_logic;
			clrn :  IN std_logic;
			ena  :  IN std_logic;
			q    : OUT std_logic_vector(3 DOWNTO 0));
END reg_pp_4bits;

ARCHITECTURE arch OF reg_pp_4bits IS
BEGIN
	PROCESS(clk, clrn)
	BEGIN
		IF(clrn='0') THEN
			q <= "0000";
		ELSIF (clk'EVENT and clk='1') THEN
			IF (ena='1') THEN
				q <= d;
			END IF;
		END IF;
	END PROCESS;
END arch;